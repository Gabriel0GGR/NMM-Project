library verilog;
use verilog.vl_types.all;
entity nmm_vlg_vec_tst is
end nmm_vlg_vec_tst;
