library verilog;
use verilog.vl_types.all;
entity NMM_vlg_vec_tst is
end NMM_vlg_vec_tst;
