library verilog;
use verilog.vl_types.all;
entity nmm_vlg_check_tst is
    port(
        c_out           : in     vl_logic;
        load            : in     vl_logic;
        pin_name1       : in     vl_logic;
        pin_name2       : in     vl_logic;
        pin_name3       : in     vl_logic;
        pin_name4       : in     vl_logic;
        pin_name5       : in     vl_logic;
        pin_name6       : in     vl_logic;
        pin_name7       : in     vl_logic;
        pin_name8       : in     vl_logic;
        pin_name9       : in     vl_logic;
        pin_name10      : in     vl_logic;
        pin_name11      : in     vl_logic;
        pin_name12      : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end nmm_vlg_check_tst;
