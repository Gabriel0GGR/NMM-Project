library verilog;
use verilog.vl_types.all;
entity clk_multiplier_vlg_vec_tst is
end clk_multiplier_vlg_vec_tst;
